// Program: 
// Author: Rajesh Kumar Bhuyan
// Date: Dec 29 2020
// Assignment: 
// Purpose: 
// 
// Input: 
// Output: 
// Related
// Files: 
// Functions: 
// 

