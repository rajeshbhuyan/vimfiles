// Program: 
// Author: Rajesh kumar Bhuyan
// Date: Dec 29 2020
// Assignment: 
// Purpose: 
// 
// Input: 
// Output: 
// Related
// Files: 
// Functions: 
// 

